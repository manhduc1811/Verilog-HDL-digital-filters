module testbench_500Hz;
    // Inputs
    reg clk, reset;
    reg signed [31:0] x;
    wire signed [31:0] y;
    // Instantiate the Unit Under Test (UUT)
    iir DUT(
      .clk(clk),
      .rst(reset),
      .x(x),
      .y(y)
    );
    // Generate clock with 100ns period
    initial clk = 0;
    always #20833 clk = ~clk;

    initial begin
        x = 32'd0;
        reset = 1;
        clk = 0;
        #10;
        reset = 0;
        #20;
        reset = 1;
        #10;
		x =                0; #20833; // Sample(1)
		x =              297; #20833; // Sample(2)
		x =             -173; #20833; // Sample(3)
		x =              -56; #20833; // Sample(4)
		x =              378; #20833; // Sample(5)
		x =              -19; #20833; // Sample(6)
		x =              -97; #20833; // Sample(7)
		x =              410; #20833; // Sample(8)
		x =              150; #20833; // Sample(9)
		x =             -110; #20833; // Sample(10)
		x =              395; #20833; // Sample(11)
		x =              313; #20833; // Sample(12)
		x =              -88; #20833; // Sample(13)
		x =              341; #20833; // Sample(14)
		x =              450; #20833; // Sample(15)
		x =              -28; #20833; // Sample(16)
		x =              260; #20833; // Sample(17)
		x =              546; #20833; // Sample(18)
		x =               65; #20833; // Sample(19)
		x =              169; #20833; // Sample(20)
		x =              590; #20833; // Sample(21)
		x =              179; #20833; // Sample(22)
		x =               85; #20833; // Sample(23)
		x =              576; #20833; // Sample(24)
		x =              300; #20833; // Sample(25)
		x =               22; #20833; // Sample(26)
		x =              509; #20833; // Sample(27)
		x =              409; #20833; // Sample(28)
		x =              -10; #20833; // Sample(29)
		x =              399; #20833; // Sample(30)
		x =              489; #20833; // Sample(31)
		x =               -8; #20833; // Sample(32)
		x =              260; #20833; // Sample(33)
		x =              526; #20833; // Sample(34)
		x =               26; #20833; // Sample(35)
		x =              111; #20833; // Sample(36)
		x =              512; #20833; // Sample(37)
		x =               83; #20833; // Sample(38)
		x =              -29; #20833; // Sample(39)
		x =              444; #20833; // Sample(40)
		x =              150; #20833; // Sample(41)
		x =             -144; #20833; // Sample(42)
		x =              327; #20833; // Sample(43)
		x =              211; #20833; // Sample(44)
		x =             -222; #20833; // Sample(45)
		x =              174; #20833; // Sample(46)
		x =              251; #20833; // Sample(47)
		x =             -257; #20833; // Sample(48)
		x =                0; #20833; // Sample(49)
		x =              257; #20833; // Sample(50)
		x =             -251; #20833; // Sample(51)
		x =             -174; #20833; // Sample(52)
		x =              222; #20833; // Sample(53)
		x =             -211; #20833; // Sample(54)
		x =             -327; #20833; // Sample(55)
		x =              144; #20833; // Sample(56)
		x =             -150; #20833; // Sample(57)
		x =             -444; #20833; // Sample(58)
		x =               29; #20833; // Sample(59)
		x =              -83; #20833; // Sample(60)
		x =             -512; #20833; // Sample(61)
		x =             -111; #20833; // Sample(62)
		x =              -26; #20833; // Sample(63)
		x =             -526; #20833; // Sample(64)
		x =             -260; #20833; // Sample(65)
		x =                8; #20833; // Sample(66)
		x =             -489; #20833; // Sample(67)
		x =             -399; #20833; // Sample(68)
		x =               10; #20833; // Sample(69)
		x =             -409; #20833; // Sample(70)
		x =             -509; #20833; // Sample(71)
		x =              -22; #20833; // Sample(72)
		x =             -300; #20833; // Sample(73)
		x =             -576; #20833; // Sample(74)
		x =              -85; #20833; // Sample(75)
		x =             -179; #20833; // Sample(76)
		x =             -590; #20833; // Sample(77)
		x =             -169; #20833; // Sample(78)
		x =              -65; #20833; // Sample(79)
		x =             -546; #20833; // Sample(80)
		x =             -260; #20833; // Sample(81)
		x =               28; #20833; // Sample(82)
		x =             -450; #20833; // Sample(83)
		x =             -341; #20833; // Sample(84)
		x =               88; #20833; // Sample(85)
		x =             -313; #20833; // Sample(86)
		x =             -395; #20833; // Sample(87)
		x =              110; #20833; // Sample(88)
		x =             -150; #20833; // Sample(89)
		x =             -410; #20833; // Sample(90)
		x =               97; #20833; // Sample(91)
		x =               19; #20833; // Sample(92)
		x =             -378; #20833; // Sample(93)
		x =               56; #20833; // Sample(94)
		x =              173; #20833; // Sample(95)
		x =             -297; #20833; // Sample(96)
		x =               -0; #20833; // Sample(97)
		x =              297; #20833; // Sample(98)
		x =             -173; #20833; // Sample(99)
		x =              -56; #20833; // Sample(100)
		x =              378; #20833; // Sample(101)
		x =              -19; #20833; // Sample(102)
		x =              -97; #20833; // Sample(103)
		x =              410; #20833; // Sample(104)
		x =              150; #20833; // Sample(105)
		x =             -110; #20833; // Sample(106)
		x =              395; #20833; // Sample(107)
		x =              313; #20833; // Sample(108)
		x =              -88; #20833; // Sample(109)
		x =              341; #20833; // Sample(110)
		x =              450; #20833; // Sample(111)
		x =              -28; #20833; // Sample(112)
		x =              260; #20833; // Sample(113)
		x =              546; #20833; // Sample(114)
		x =               65; #20833; // Sample(115)
		x =              169; #20833; // Sample(116)
		x =              590; #20833; // Sample(117)
		x =              179; #20833; // Sample(118)
		x =               85; #20833; // Sample(119)
		x =              576; #20833; // Sample(120)
		x =              300; #20833; // Sample(121)
		x =               22; #20833; // Sample(122)
		x =              509; #20833; // Sample(123)
		x =              409; #20833; // Sample(124)
		x =              -10; #20833; // Sample(125)
		x =              399; #20833; // Sample(126)
		x =              489; #20833; // Sample(127)
		x =               -8; #20833; // Sample(128)
		x =              260; #20833; // Sample(129)
		x =              526; #20833; // Sample(130)
		x =               26; #20833; // Sample(131)
		x =              111; #20833; // Sample(132)
		x =              512; #20833; // Sample(133)
		x =               83; #20833; // Sample(134)
		x =              -29; #20833; // Sample(135)
		x =              444; #20833; // Sample(136)
		x =              150; #20833; // Sample(137)
		x =             -144; #20833; // Sample(138)
		x =              327; #20833; // Sample(139)
		x =              211; #20833; // Sample(140)
		x =             -222; #20833; // Sample(141)
		x =              174; #20833; // Sample(142)
		x =              251; #20833; // Sample(143)
		x =             -257; #20833; // Sample(144)
		x =                0; #20833; // Sample(145)
		x =              257; #20833; // Sample(146)
		x =             -251; #20833; // Sample(147)
		x =             -174; #20833; // Sample(148)
		x =              222; #20833; // Sample(149)
		x =             -211; #20833; // Sample(150)
		x =             -327; #20833; // Sample(151)
		x =              144; #20833; // Sample(152)
		x =             -150; #20833; // Sample(153)
		x =             -444; #20833; // Sample(154)
		x =               29; #20833; // Sample(155)
		x =              -83; #20833; // Sample(156)
		x =             -512; #20833; // Sample(157)
		x =             -111; #20833; // Sample(158)
		x =              -26; #20833; // Sample(159)
		x =             -526; #20833; // Sample(160)
		x =             -260; #20833; // Sample(161)
		x =                8; #20833; // Sample(162)
		x =             -489; #20833; // Sample(163)
		x =             -399; #20833; // Sample(164)
		x =               10; #20833; // Sample(165)
		x =             -409; #20833; // Sample(166)
		x =             -509; #20833; // Sample(167)
		x =              -22; #20833; // Sample(168)
		x =             -300; #20833; // Sample(169)
		x =             -576; #20833; // Sample(170)
		x =              -85; #20833; // Sample(171)
		x =             -179; #20833; // Sample(172)
		x =             -590; #20833; // Sample(173)
		x =             -169; #20833; // Sample(174)
		x =              -65; #20833; // Sample(175)
		x =             -546; #20833; // Sample(176)
		x =             -260; #20833; // Sample(177)
		x =               28; #20833; // Sample(178)
		x =             -450; #20833; // Sample(179)
		x =             -341; #20833; // Sample(180)
		x =               88; #20833; // Sample(181)
		x =             -313; #20833; // Sample(182)
		x =             -395; #20833; // Sample(183)
		x =              110; #20833; // Sample(184)
		x =             -150; #20833; // Sample(185)
		x =             -410; #20833; // Sample(186)
		x =               97; #20833; // Sample(187)
		x =               19; #20833; // Sample(188)
		x =             -378; #20833; // Sample(189)
		x =               56; #20833; // Sample(190)
		x =              173; #20833; // Sample(191)
		x =             -297; #20833; // Sample(192)
		x =               -0; #20833; // Sample(193)
		x =              297; #20833; // Sample(194)
		x =             -173; #20833; // Sample(195)
		x =              -56; #20833; // Sample(196)
		x =              378; #20833; // Sample(197)
		x =              -19; #20833; // Sample(198)
		x =              -97; #20833; // Sample(199)
		x =              410; #20833; // Sample(200)
		x =              150; #20833; // Sample(201)
		x =             -110; #20833; // Sample(202)
		x =              395; #20833; // Sample(203)
		x =              313; #20833; // Sample(204)
		x =              -88; #20833; // Sample(205)
		x =              341; #20833; // Sample(206)
		x =              450; #20833; // Sample(207)
		x =              -28; #20833; // Sample(208)
		x =              260; #20833; // Sample(209)
		x =              546; #20833; // Sample(210)
		x =               65; #20833; // Sample(211)
		x =              169; #20833; // Sample(212)
		x =              590; #20833; // Sample(213)
		x =              179; #20833; // Sample(214)
		x =               85; #20833; // Sample(215)
		x =              576; #20833; // Sample(216)
		x =              300; #20833; // Sample(217)
		x =               22; #20833; // Sample(218)
		x =              509; #20833; // Sample(219)
		x =              409; #20833; // Sample(220)
		x =              -10; #20833; // Sample(221)
		x =              399; #20833; // Sample(222)
		x =              489; #20833; // Sample(223)
		x =               -8; #20833; // Sample(224)
		x =              260; #20833; // Sample(225)
		x =              526; #20833; // Sample(226)
		x =               26; #20833; // Sample(227)
		x =              111; #20833; // Sample(228)
		x =              512; #20833; // Sample(229)
		x =               83; #20833; // Sample(230)
		x =              -29; #20833; // Sample(231)
		x =              444; #20833; // Sample(232)
		x =              150; #20833; // Sample(233)
		x =             -144; #20833; // Sample(234)
		x =              327; #20833; // Sample(235)
		x =              211; #20833; // Sample(236)
		x =             -222; #20833; // Sample(237)
		x =              174; #20833; // Sample(238)
		x =              251; #20833; // Sample(239)
		x =             -257; #20833; // Sample(240)
		x =                0; #20833; // Sample(241)
		x =              257; #20833; // Sample(242)
		x =             -251; #20833; // Sample(243)
		x =             -174; #20833; // Sample(244)
		x =              222; #20833; // Sample(245)
		x =             -211; #20833; // Sample(246)
		x =             -327; #20833; // Sample(247)
		x =              144; #20833; // Sample(248)
		x =             -150; #20833; // Sample(249)
		x =             -444; #20833; // Sample(250)
		x =               29; #20833; // Sample(251)
		x =              -83; #20833; // Sample(252)
		x =             -512; #20833; // Sample(253)
		x =             -111; #20833; // Sample(254)
		x =              -26; #20833; // Sample(255)
		x =             -526; #20833; // Sample(256)
		x =             -260; #20833; // Sample(257)
		x =                8; #20833; // Sample(258)
		x =             -489; #20833; // Sample(259)
		x =             -399; #20833; // Sample(260)
		x =               10; #20833; // Sample(261)
		x =             -409; #20833; // Sample(262)
		x =             -509; #20833; // Sample(263)
		x =              -22; #20833; // Sample(264)
		x =             -300; #20833; // Sample(265)
		x =             -576; #20833; // Sample(266)
		x =              -85; #20833; // Sample(267)
		x =             -179; #20833; // Sample(268)
		x =             -590; #20833; // Sample(269)
		x =             -169; #20833; // Sample(270)
		x =              -65; #20833; // Sample(271)
		x =             -546; #20833; // Sample(272)
		x =             -260; #20833; // Sample(273)
		x =               28; #20833; // Sample(274)
		x =             -450; #20833; // Sample(275)
		x =             -341; #20833; // Sample(276)
		x =               88; #20833; // Sample(277)
		x =             -313; #20833; // Sample(278)
		x =             -395; #20833; // Sample(279)
		x =              110; #20833; // Sample(280)
		x =             -150; #20833; // Sample(281)
		x =             -410; #20833; // Sample(282)
		x =               97; #20833; // Sample(283)
		x =               19; #20833; // Sample(284)
		x =             -378; #20833; // Sample(285)
		x =               56; #20833; // Sample(286)
		x =              173; #20833; // Sample(287)
		x =             -297; #20833; // Sample(288)
		x =               -0; #20833; // Sample(289)
		x =              297; #20833; // Sample(290)
		x =             -173; #20833; // Sample(291)
		x =              -56; #20833; // Sample(292)
		x =              378; #20833; // Sample(293)
		x =              -19; #20833; // Sample(294)
		x =              -97; #20833; // Sample(295)
		x =              410; #20833; // Sample(296)
		x =              150; #20833; // Sample(297)
		x =             -110; #20833; // Sample(298)
		x =              395; #20833; // Sample(299)
		x =              313; #20833; // Sample(300)
		x =              -88; #20833; // Sample(301)
		x =              341; #20833; // Sample(302)
		x =              450; #20833; // Sample(303)
		x =              -28; #20833; // Sample(304)
		x =              260; #20833; // Sample(305)
		x =              546; #20833; // Sample(306)
		x =               65; #20833; // Sample(307)
		x =              169; #20833; // Sample(308)
		x =              590; #20833; // Sample(309)
		x =              179; #20833; // Sample(310)
		x =               85; #20833; // Sample(311)
		x =              576; #20833; // Sample(312)
		x =              300; #20833; // Sample(313)
		x =               22; #20833; // Sample(314)
		x =              509; #20833; // Sample(315)
		x =              409; #20833; // Sample(316)
		x =              -10; #20833; // Sample(317)
		x =              399; #20833; // Sample(318)
		x =              489; #20833; // Sample(319)
		x =               -8; #20833; // Sample(320)
		x =              260; #20833; // Sample(321)
		x =              526; #20833; // Sample(322)
		x =               26; #20833; // Sample(323)
		x =              111; #20833; // Sample(324)
		x =              512; #20833; // Sample(325)
		x =               83; #20833; // Sample(326)
		x =              -29; #20833; // Sample(327)
		x =              444; #20833; // Sample(328)
		x =              150; #20833; // Sample(329)
		x =             -144; #20833; // Sample(330)
		x =              327; #20833; // Sample(331)
		x =              211; #20833; // Sample(332)
		x =             -222; #20833; // Sample(333)
		x =              174; #20833; // Sample(334)
		x =              251; #20833; // Sample(335)
		x =             -257; #20833; // Sample(336)
		x =                0; #20833; // Sample(337)
		x =              257; #20833; // Sample(338)
		x =             -251; #20833; // Sample(339)
		x =             -174; #20833; // Sample(340)
		x =              222; #20833; // Sample(341)
		x =             -211; #20833; // Sample(342)
		x =             -327; #20833; // Sample(343)
		x =              144; #20833; // Sample(344)
		x =             -150; #20833; // Sample(345)
		x =             -444; #20833; // Sample(346)
		x =               29; #20833; // Sample(347)
		x =              -83; #20833; // Sample(348)
		x =             -512; #20833; // Sample(349)
		x =             -111; #20833; // Sample(350)
		x =              -26; #20833; // Sample(351)
		x =             -526; #20833; // Sample(352)
		x =             -260; #20833; // Sample(353)
		x =                8; #20833; // Sample(354)
		x =             -489; #20833; // Sample(355)
		x =             -399; #20833; // Sample(356)
		x =               10; #20833; // Sample(357)
		x =             -409; #20833; // Sample(358)
		x =             -509; #20833; // Sample(359)
		x =              -22; #20833; // Sample(360)
		x =             -300; #20833; // Sample(361)
		x =             -576; #20833; // Sample(362)
		x =              -85; #20833; // Sample(363)
		x =             -179; #20833; // Sample(364)
		x =             -590; #20833; // Sample(365)
		x =             -169; #20833; // Sample(366)
		x =              -65; #20833; // Sample(367)
		x =             -546; #20833; // Sample(368)
		x =             -260; #20833; // Sample(369)
		x =               28; #20833; // Sample(370)
		x =             -450; #20833; // Sample(371)
		x =             -341; #20833; // Sample(372)
		x =               88; #20833; // Sample(373)
		x =             -313; #20833; // Sample(374)
		x =             -395; #20833; // Sample(375)
		x =              110; #20833; // Sample(376)
		x =             -150; #20833; // Sample(377)
		x =             -410; #20833; // Sample(378)
		x =               97; #20833; // Sample(379)
		x =               19; #20833; // Sample(380)
		x =             -378; #20833; // Sample(381)
		x =               56; #20833; // Sample(382)
		x =              173; #20833; // Sample(383)
		x =             -297; #20833; // Sample(384)
		x =               -0; #20833; // Sample(385)
		x =              297; #20833; // Sample(386)
		x =             -173; #20833; // Sample(387)
		x =              -56; #20833; // Sample(388)
		x =              378; #20833; // Sample(389)
		x =              -19; #20833; // Sample(390)
		x =              -97; #20833; // Sample(391)
		x =              410; #20833; // Sample(392)
		x =              150; #20833; // Sample(393)
		x =             -110; #20833; // Sample(394)
		x =              395; #20833; // Sample(395)
		x =              313; #20833; // Sample(396)
		x =              -88; #20833; // Sample(397)
		x =              341; #20833; // Sample(398)
		x =              450; #20833; // Sample(399)
		x =              -28; #20833; // Sample(400)
		x =              260; #20833; // Sample(401)
		x =              546; #20833; // Sample(402)
		x =               65; #20833; // Sample(403)
		x =              169; #20833; // Sample(404)
		x =              590; #20833; // Sample(405)
		x =              179; #20833; // Sample(406)
		x =               85; #20833; // Sample(407)
		x =              576; #20833; // Sample(408)
		x =              300; #20833; // Sample(409)
		x =               22; #20833; // Sample(410)
		x =              509; #20833; // Sample(411)
		x =              409; #20833; // Sample(412)
		x =              -10; #20833; // Sample(413)
		x =              399; #20833; // Sample(414)
		x =              489; #20833; // Sample(415)
		x =               -8; #20833; // Sample(416)
		x =              260; #20833; // Sample(417)
		x =              526; #20833; // Sample(418)
		x =               26; #20833; // Sample(419)
		x =              111; #20833; // Sample(420)
		x =              512; #20833; // Sample(421)
		x =               83; #20833; // Sample(422)
		x =              -29; #20833; // Sample(423)
		x =              444; #20833; // Sample(424)
		x =              150; #20833; // Sample(425)
		x =             -144; #20833; // Sample(426)
		x =              327; #20833; // Sample(427)
		x =              211; #20833; // Sample(428)
		x =             -222; #20833; // Sample(429)
		x =              174; #20833; // Sample(430)
		x =              251; #20833; // Sample(431)
		x =             -257; #20833; // Sample(432)
		x =                0; #20833; // Sample(433)
		x =              257; #20833; // Sample(434)
		x =             -251; #20833; // Sample(435)
		x =             -174; #20833; // Sample(436)
		x =              222; #20833; // Sample(437)
		x =             -211; #20833; // Sample(438)
		x =             -327; #20833; // Sample(439)
		x =              144; #20833; // Sample(440)
		x =             -150; #20833; // Sample(441)
		x =             -444; #20833; // Sample(442)
		x =               29; #20833; // Sample(443)
		x =              -83; #20833; // Sample(444)
		x =             -512; #20833; // Sample(445)
		x =             -111; #20833; // Sample(446)
		x =              -26; #20833; // Sample(447)
		x =             -526; #20833; // Sample(448)
		x =             -260; #20833; // Sample(449)
		x =                8; #20833; // Sample(450)
		x =             -489; #20833; // Sample(451)
		x =             -399; #20833; // Sample(452)
		x =               10; #20833; // Sample(453)
		x =             -409; #20833; // Sample(454)
		x =             -509; #20833; // Sample(455)
		x =              -22; #20833; // Sample(456)
		x =             -300; #20833; // Sample(457)
		x =             -576; #20833; // Sample(458)
		x =              -85; #20833; // Sample(459)
		x =             -179; #20833; // Sample(460)
		x =             -590; #20833; // Sample(461)
		x =             -169; #20833; // Sample(462)
		x =              -65; #20833; // Sample(463)
		x =             -546; #20833; // Sample(464)
		x =             -260; #20833; // Sample(465)
		x =               28; #20833; // Sample(466)
		x =             -450; #20833; // Sample(467)
		x =             -341; #20833; // Sample(468)
		x =               88; #20833; // Sample(469)
		x =             -313; #20833; // Sample(470)
		x =             -395; #20833; // Sample(471)
		x =              110; #20833; // Sample(472)
		x =             -150; #20833; // Sample(473)
		x =             -410; #20833; // Sample(474)
		x =               97; #20833; // Sample(475)
		x =               19; #20833; // Sample(476)
		x =             -378; #20833; // Sample(477)
		x =               56; #20833; // Sample(478)
		x =              173; #20833; // Sample(479)
		x =             -297; #20833; // Sample(480)
		x =               -0; #20833; // Sample(481)
		x =              297; #20833; // Sample(482)
		x =             -173; #20833; // Sample(483)
		x =              -56; #20833; // Sample(484)
		x =              378; #20833; // Sample(485)
		x =              -19; #20833; // Sample(486)
		x =              -97; #20833; // Sample(487)
		x =              410; #20833; // Sample(488)
		x =              150; #20833; // Sample(489)
		x =             -110; #20833; // Sample(490)
		x =              395; #20833; // Sample(491)
		x =              313; #20833; // Sample(492)
		x =              -88; #20833; // Sample(493)
		x =              341; #20833; // Sample(494)
		x =              450; #20833; // Sample(495)
		x =              -28; #20833; // Sample(496)
		x =              260; #20833; // Sample(497)
		x =              546; #20833; // Sample(498)
		x =               65; #20833; // Sample(499)
		x =              169; #20833; // Sample(500)
		x =                0; #20833; // Sample(501)
		x =              183; #20833; // Sample(502)
		x =              290; #20833; // Sample(503)
		x =              277; #20833; // Sample(504)
		x =              150; #20833; // Sample(505)
		x =              -39; #20833; // Sample(506)
		x =             -212; #20833; // Sample(507)
		x =             -297; #20833; // Sample(508)
		x =             -260; #20833; // Sample(509)
		x =             -115; #20833; // Sample(510)
		x =               78; #20833; // Sample(511)
		x =              238; #20833; // Sample(512)
		x =              300; #20833; // Sample(513)
		x =              238; #20833; // Sample(514)
		x =               78; #20833; // Sample(515)
		x =             -115; #20833; // Sample(516)
		x =             -260; #20833; // Sample(517)
		x =             -297; #20833; // Sample(518)
		x =             -212; #20833; // Sample(519)
		x =              -39; #20833; // Sample(520)
		x =              150; #20833; // Sample(521)
		x =              277; #20833; // Sample(522)
		x =              290; #20833; // Sample(523)
		x =              183; #20833; // Sample(524)
		x =                0; #20833; // Sample(525)
		x =             -183; #20833; // Sample(526)
		x =             -290; #20833; // Sample(527)
		x =             -277; #20833; // Sample(528)
		x =             -150; #20833; // Sample(529)
		x =               39; #20833; // Sample(530)
		x =              212; #20833; // Sample(531)
		x =              297; #20833; // Sample(532)
		x =              260; #20833; // Sample(533)
		x =              115; #20833; // Sample(534)
		x =              -78; #20833; // Sample(535)
		x =             -238; #20833; // Sample(536)
		x =             -300; #20833; // Sample(537)
		x =             -238; #20833; // Sample(538)
		x =              -78; #20833; // Sample(539)
		x =              115; #20833; // Sample(540)
		x =              260; #20833; // Sample(541)
		x =              297; #20833; // Sample(542)
		x =              212; #20833; // Sample(543)
		x =               39; #20833; // Sample(544)
		x =             -150; #20833; // Sample(545)
		x =             -277; #20833; // Sample(546)
		x =             -290; #20833; // Sample(547)
		x =             -183; #20833; // Sample(548)
		x =               -0; #20833; // Sample(549)
		x =              183; #20833; // Sample(550)
		x =              290; #20833; // Sample(551)
		x =              277; #20833; // Sample(552)
		x =              150; #20833; // Sample(553)
		x =              -39; #20833; // Sample(554)
		x =             -212; #20833; // Sample(555)
		x =             -297; #20833; // Sample(556)
		x =             -260; #20833; // Sample(557)
		x =             -115; #20833; // Sample(558)
		x =               78; #20833; // Sample(559)
		x =              238; #20833; // Sample(560)
		x =              300; #20833; // Sample(561)
		x =              238; #20833; // Sample(562)
		x =               78; #20833; // Sample(563)
		x =             -115; #20833; // Sample(564)
		x =             -260; #20833; // Sample(565)
		x =             -297; #20833; // Sample(566)
		x =             -212; #20833; // Sample(567)
		x =              -39; #20833; // Sample(568)
		x =              150; #20833; // Sample(569)
		x =              277; #20833; // Sample(570)
		x =              290; #20833; // Sample(571)
		x =              183; #20833; // Sample(572)
		x =               -0; #20833; // Sample(573)
		x =             -183; #20833; // Sample(574)
		x =             -290; #20833; // Sample(575)
		x =             -277; #20833; // Sample(576)
		x =             -150; #20833; // Sample(577)
		x =               39; #20833; // Sample(578)
		x =              212; #20833; // Sample(579)
		x =              297; #20833; // Sample(580)
		x =              260; #20833; // Sample(581)
		x =              115; #20833; // Sample(582)
		x =              -78; #20833; // Sample(583)
		x =             -238; #20833; // Sample(584)
		x =             -300; #20833; // Sample(585)
		x =             -238; #20833; // Sample(586)
		x =              -78; #20833; // Sample(587)
		x =              115; #20833; // Sample(588)
		x =              260; #20833; // Sample(589)
		x =              297; #20833; // Sample(590)
		x =              212; #20833; // Sample(591)
		x =               39; #20833; // Sample(592)
		x =             -150; #20833; // Sample(593)
		x =             -277; #20833; // Sample(594)
		x =             -290; #20833; // Sample(595)
		x =             -183; #20833; // Sample(596)
		x =               -0; #20833; // Sample(597)
		x =              183; #20833; // Sample(598)
		x =              290; #20833; // Sample(599)
		x =              277; #20833; // Sample(600)
		x =              150; #20833; // Sample(601)
		x =              -39; #20833; // Sample(602)
		x =             -212; #20833; // Sample(603)
		x =             -297; #20833; // Sample(604)
		x =             -260; #20833; // Sample(605)
		x =             -115; #20833; // Sample(606)
		x =               78; #20833; // Sample(607)
		x =              238; #20833; // Sample(608)
		x =              300; #20833; // Sample(609)
		x =              238; #20833; // Sample(610)
		x =               78; #20833; // Sample(611)
		x =             -115; #20833; // Sample(612)
		x =             -260; #20833; // Sample(613)
		x =             -297; #20833; // Sample(614)
		x =             -212; #20833; // Sample(615)
		x =              -39; #20833; // Sample(616)
		x =              150; #20833; // Sample(617)
		x =              277; #20833; // Sample(618)
		x =              290; #20833; // Sample(619)
		x =              183; #20833; // Sample(620)
		x =               -0; #20833; // Sample(621)
		x =             -183; #20833; // Sample(622)
		x =             -290; #20833; // Sample(623)
		x =             -277; #20833; // Sample(624)
		x =             -150; #20833; // Sample(625)
		x =               39; #20833; // Sample(626)
		x =              212; #20833; // Sample(627)
		x =              297; #20833; // Sample(628)
		x =              260; #20833; // Sample(629)
		x =              115; #20833; // Sample(630)
		x =              -78; #20833; // Sample(631)
		x =             -238; #20833; // Sample(632)
		x =             -300; #20833; // Sample(633)
		x =             -238; #20833; // Sample(634)
		x =              -78; #20833; // Sample(635)
		x =              115; #20833; // Sample(636)
		x =              260; #20833; // Sample(637)
		x =              297; #20833; // Sample(638)
		x =              212; #20833; // Sample(639)
		x =               39; #20833; // Sample(640)
		x =             -150; #20833; // Sample(641)
		x =             -277; #20833; // Sample(642)
		x =             -290; #20833; // Sample(643)
		x =             -183; #20833; // Sample(644)
		x =                0; #20833; // Sample(645)
		x =              183; #20833; // Sample(646)
		x =              290; #20833; // Sample(647)
		x =              277; #20833; // Sample(648)
		x =              150; #20833; // Sample(649)
		x =              -39; #20833; // Sample(650)
		x =             -212; #20833; // Sample(651)
		x =             -297; #20833; // Sample(652)
		x =             -260; #20833; // Sample(653)
		x =             -115; #20833; // Sample(654)
		x =               78; #20833; // Sample(655)
		x =              238; #20833; // Sample(656)
		x =              300; #20833; // Sample(657)
		x =              238; #20833; // Sample(658)
		x =               78; #20833; // Sample(659)
		x =             -115; #20833; // Sample(660)
		x =             -260; #20833; // Sample(661)
		x =             -297; #20833; // Sample(662)
		x =             -212; #20833; // Sample(663)
		x =              -39; #20833; // Sample(664)
		x =              150; #20833; // Sample(665)
		x =              277; #20833; // Sample(666)
		x =              290; #20833; // Sample(667)
		x =              183; #20833; // Sample(668)
		x =               -0; #20833; // Sample(669)
		x =             -183; #20833; // Sample(670)
		x =             -290; #20833; // Sample(671)
		x =             -277; #20833; // Sample(672)
		x =             -150; #20833; // Sample(673)
		x =               39; #20833; // Sample(674)
		x =              212; #20833; // Sample(675)
		x =              297; #20833; // Sample(676)
		x =              260; #20833; // Sample(677)
		x =              115; #20833; // Sample(678)
		x =              -78; #20833; // Sample(679)
		x =             -238; #20833; // Sample(680)
		x =             -300; #20833; // Sample(681)
		x =             -238; #20833; // Sample(682)
		x =              -78; #20833; // Sample(683)
		x =              115; #20833; // Sample(684)
		x =              260; #20833; // Sample(685)
		x =              297; #20833; // Sample(686)
		x =              212; #20833; // Sample(687)
		x =               39; #20833; // Sample(688)
		x =             -150; #20833; // Sample(689)
		x =             -277; #20833; // Sample(690)
		x =             -290; #20833; // Sample(691)
		x =             -183; #20833; // Sample(692)
		x =               -0; #20833; // Sample(693)
		x =              183; #20833; // Sample(694)
		x =              290; #20833; // Sample(695)
		x =              277; #20833; // Sample(696)
		x =              150; #20833; // Sample(697)
		x =              -39; #20833; // Sample(698)
		x =             -212; #20833; // Sample(699)
		x =             -297; #20833; // Sample(700)
		x =             -260; #20833; // Sample(701)
		x =             -115; #20833; // Sample(702)
		x =               78; #20833; // Sample(703)
		x =              238; #20833; // Sample(704)
		x =              300; #20833; // Sample(705)
		x =              238; #20833; // Sample(706)
		x =               78; #20833; // Sample(707)
		x =             -115; #20833; // Sample(708)
		x =             -260; #20833; // Sample(709)
		x =             -297; #20833; // Sample(710)
		x =             -212; #20833; // Sample(711)
		x =              -39; #20833; // Sample(712)
		x =              150; #20833; // Sample(713)
		x =              277; #20833; // Sample(714)
		x =              290; #20833; // Sample(715)
		x =              183; #20833; // Sample(716)
		x =                0; #20833; // Sample(717)
		x =             -183; #20833; // Sample(718)
		x =             -290; #20833; // Sample(719)
		x =             -277; #20833; // Sample(720)
		x =             -150; #20833; // Sample(721)
		x =               39; #20833; // Sample(722)
		x =              212; #20833; // Sample(723)
		x =              297; #20833; // Sample(724)
		x =              260; #20833; // Sample(725)
		x =              115; #20833; // Sample(726)
		x =              -78; #20833; // Sample(727)
		x =             -238; #20833; // Sample(728)
		x =             -300; #20833; // Sample(729)
		x =             -238; #20833; // Sample(730)
		x =              -78; #20833; // Sample(731)
		x =              115; #20833; // Sample(732)
		x =              260; #20833; // Sample(733)
		x =              297; #20833; // Sample(734)
		x =              212; #20833; // Sample(735)
		x =               39; #20833; // Sample(736)
		x =             -150; #20833; // Sample(737)
		x =             -277; #20833; // Sample(738)
		x =             -290; #20833; // Sample(739)
		x =             -183; #20833; // Sample(740)
		x =                0; #20833; // Sample(741)
		x =              183; #20833; // Sample(742)
		x =              290; #20833; // Sample(743)
		x =              277; #20833; // Sample(744)
		x =              150; #20833; // Sample(745)
		x =              -39; #20833; // Sample(746)
		x =             -212; #20833; // Sample(747)
		x =             -297; #20833; // Sample(748)
		x =             -260; #20833; // Sample(749)
		x =             -115; #20833; // Sample(750)
		x =               78; #20833; // Sample(751)
		x =              238; #20833; // Sample(752)
		x =              300; #20833; // Sample(753)
		x =              238; #20833; // Sample(754)
		x =               78; #20833; // Sample(755)
		x =             -115; #20833; // Sample(756)
		x =             -260; #20833; // Sample(757)
		x =             -297; #20833; // Sample(758)
		x =             -212; #20833; // Sample(759)
		x =              -39; #20833; // Sample(760)
		x =              150; #20833; // Sample(761)
		x =              277; #20833; // Sample(762)
		x =              290; #20833; // Sample(763)
		x =              183; #20833; // Sample(764)
		x =               -0; #20833; // Sample(765)
		x =             -183; #20833; // Sample(766)
		x =             -290; #20833; // Sample(767)
		x =             -277; #20833; // Sample(768)
		x =             -150; #20833; // Sample(769)
		x =               39; #20833; // Sample(770)
		x =              212; #20833; // Sample(771)
		x =              297; #20833; // Sample(772)
		x =              260; #20833; // Sample(773)
		x =              115; #20833; // Sample(774)
		x =              -78; #20833; // Sample(775)
		x =             -238; #20833; // Sample(776)
		x =             -300; #20833; // Sample(777)
		x =             -238; #20833; // Sample(778)
		x =              -78; #20833; // Sample(779)
		x =              115; #20833; // Sample(780)
		x =              260; #20833; // Sample(781)
		x =              297; #20833; // Sample(782)
		x =              212; #20833; // Sample(783)
		x =               39; #20833; // Sample(784)
		x =             -150; #20833; // Sample(785)
		x =             -277; #20833; // Sample(786)
		x =             -290; #20833; // Sample(787)
		x =             -183; #20833; // Sample(788)
		x =                0; #20833; // Sample(789)
		x =              183; #20833; // Sample(790)
		x =              290; #20833; // Sample(791)
		x =              277; #20833; // Sample(792)
		x =              150; #20833; // Sample(793)
		x =              -39; #20833; // Sample(794)
		x =             -212; #20833; // Sample(795)
		x =             -297; #20833; // Sample(796)
		x =             -260; #20833; // Sample(797)
		x =             -115; #20833; // Sample(798)
		x =               78; #20833; // Sample(799)
		x =              238; #20833; // Sample(800)
		x =              300; #20833; // Sample(801)
		x =              238; #20833; // Sample(802)
		x =               78; #20833; // Sample(803)
		x =             -115; #20833; // Sample(804)
		x =             -260; #20833; // Sample(805)
		x =             -297; #20833; // Sample(806)
		x =             -212; #20833; // Sample(807)
		x =              -39; #20833; // Sample(808)
		x =              150; #20833; // Sample(809)
		x =              277; #20833; // Sample(810)
		x =              290; #20833; // Sample(811)
		x =              183; #20833; // Sample(812)
		x =               -0; #20833; // Sample(813)
		x =             -183; #20833; // Sample(814)
		x =             -290; #20833; // Sample(815)
		x =             -277; #20833; // Sample(816)
		x =             -150; #20833; // Sample(817)
		x =               39; #20833; // Sample(818)
		x =              212; #20833; // Sample(819)
		x =              297; #20833; // Sample(820)
		x =              260; #20833; // Sample(821)
		x =              115; #20833; // Sample(822)
		x =              -78; #20833; // Sample(823)
		x =             -238; #20833; // Sample(824)
		x =             -300; #20833; // Sample(825)
		x =             -238; #20833; // Sample(826)
		x =              -78; #20833; // Sample(827)
		x =              115; #20833; // Sample(828)
		x =              260; #20833; // Sample(829)
		x =              297; #20833; // Sample(830)
		x =              212; #20833; // Sample(831)
		x =               39; #20833; // Sample(832)
		x =             -150; #20833; // Sample(833)
		x =             -277; #20833; // Sample(834)
		x =             -290; #20833; // Sample(835)
		x =             -183; #20833; // Sample(836)
		x =                0; #20833; // Sample(837)
		x =              183; #20833; // Sample(838)
		x =              290; #20833; // Sample(839)
		x =              277; #20833; // Sample(840)
		x =              150; #20833; // Sample(841)
		x =              -39; #20833; // Sample(842)
		x =             -212; #20833; // Sample(843)
		x =             -297; #20833; // Sample(844)
		x =             -260; #20833; // Sample(845)
		x =             -115; #20833; // Sample(846)
		x =               78; #20833; // Sample(847)
		x =              238; #20833; // Sample(848)
		x =              300; #20833; // Sample(849)
		x =              238; #20833; // Sample(850)
		x =               78; #20833; // Sample(851)
		x =             -115; #20833; // Sample(852)
		x =             -260; #20833; // Sample(853)
		x =             -297; #20833; // Sample(854)
		x =             -212; #20833; // Sample(855)
		x =              -39; #20833; // Sample(856)
		x =              150; #20833; // Sample(857)
		x =              277; #20833; // Sample(858)
		x =              290; #20833; // Sample(859)
		x =              183; #20833; // Sample(860)
		x =               -0; #20833; // Sample(861)
		x =             -183; #20833; // Sample(862)
		x =             -290; #20833; // Sample(863)
		x =             -277; #20833; // Sample(864)
		x =             -150; #20833; // Sample(865)
		x =               39; #20833; // Sample(866)
		x =              212; #20833; // Sample(867)
		x =              297; #20833; // Sample(868)
		x =              260; #20833; // Sample(869)
		x =              115; #20833; // Sample(870)
		x =              -78; #20833; // Sample(871)
		x =             -238; #20833; // Sample(872)
		x =             -300; #20833; // Sample(873)
		x =             -238; #20833; // Sample(874)
		x =              -78; #20833; // Sample(875)
		x =              115; #20833; // Sample(876)
		x =              260; #20833; // Sample(877)
		x =              297; #20833; // Sample(878)
		x =              212; #20833; // Sample(879)
		x =               39; #20833; // Sample(880)
		x =             -150; #20833; // Sample(881)
		x =             -277; #20833; // Sample(882)
		x =             -290; #20833; // Sample(883)
		x =             -183; #20833; // Sample(884)
		x =               -0; #20833; // Sample(885)
		x =              183; #20833; // Sample(886)
		x =              290; #20833; // Sample(887)
		x =              277; #20833; // Sample(888)
		x =              150; #20833; // Sample(889)
		x =              -39; #20833; // Sample(890)
		x =             -212; #20833; // Sample(891)
		x =             -297; #20833; // Sample(892)
		x =             -260; #20833; // Sample(893)
		x =             -115; #20833; // Sample(894)
		x =               78; #20833; // Sample(895)
		x =              238; #20833; // Sample(896)
		x =              300; #20833; // Sample(897)
		x =              238; #20833; // Sample(898)
		x =               78; #20833; // Sample(899)
		x =             -115; #20833; // Sample(900)
		x =             -260; #20833; // Sample(901)
		x =             -297; #20833; // Sample(902)
		x =             -212; #20833; // Sample(903)
		x =              -39; #20833; // Sample(904)
		x =              150; #20833; // Sample(905)
		x =              277; #20833; // Sample(906)
		x =              290; #20833; // Sample(907)
		x =              183; #20833; // Sample(908)
		x =                0; #20833; // Sample(909)
		x =             -183; #20833; // Sample(910)
		x =             -290; #20833; // Sample(911)
		x =             -277; #20833; // Sample(912)
		x =             -150; #20833; // Sample(913)
		x =               39; #20833; // Sample(914)
		x =              212; #20833; // Sample(915)
		x =              297; #20833; // Sample(916)
		x =              260; #20833; // Sample(917)
		x =              115; #20833; // Sample(918)
		x =              -78; #20833; // Sample(919)
		x =             -238; #20833; // Sample(920)
		x =             -300; #20833; // Sample(921)
		x =             -238; #20833; // Sample(922)
		x =              -78; #20833; // Sample(923)
		x =              115; #20833; // Sample(924)
		x =              260; #20833; // Sample(925)
		x =              297; #20833; // Sample(926)
		x =              212; #20833; // Sample(927)
		x =               39; #20833; // Sample(928)
		x =             -150; #20833; // Sample(929)
		x =             -277; #20833; // Sample(930)
		x =             -290; #20833; // Sample(931)
		x =             -183; #20833; // Sample(932)
		x =               -0; #20833; // Sample(933)
		x =              183; #20833; // Sample(934)
		x =              290; #20833; // Sample(935)
		x =              277; #20833; // Sample(936)
		x =              150; #20833; // Sample(937)
		x =              -39; #20833; // Sample(938)
		x =             -212; #20833; // Sample(939)
		x =             -297; #20833; // Sample(940)
		x =             -260; #20833; // Sample(941)
		x =             -115; #20833; // Sample(942)
		x =               78; #20833; // Sample(943)
		x =              238; #20833; // Sample(944)
		x =              300; #20833; // Sample(945)
		x =              238; #20833; // Sample(946)
		x =               78; #20833; // Sample(947)
		x =             -115; #20833; // Sample(948)
		x =             -260; #20833; // Sample(949)
		x =             -297; #20833; // Sample(950)
		x =             -212; #20833; // Sample(951)
		x =              -39; #20833; // Sample(952)
		x =              150; #20833; // Sample(953)
		x =              277; #20833; // Sample(954)
		x =              290; #20833; // Sample(955)
		x =              183; #20833; // Sample(956)
		x =                0; #20833; // Sample(957)
		x =             -183; #20833; // Sample(958)
		x =             -290; #20833; // Sample(959)
		x =             -277; #20833; // Sample(960)
		x =             -150; #20833; // Sample(961)
		x =               39; #20833; // Sample(962)
		x =              212; #20833; // Sample(963)
		x =              297; #20833; // Sample(964)
		x =              260; #20833; // Sample(965)
		x =              115; #20833; // Sample(966)
		x =              -78; #20833; // Sample(967)
		x =             -238; #20833; // Sample(968)
		x =             -300; #20833; // Sample(969)
		x =             -238; #20833; // Sample(970)
		x =              -78; #20833; // Sample(971)
		x =              115; #20833; // Sample(972)
		x =              260; #20833; // Sample(973)
		x =              297; #20833; // Sample(974)
		x =              212; #20833; // Sample(975)
		x =               39; #20833; // Sample(976)
		x =             -150; #20833; // Sample(977)
		x =             -277; #20833; // Sample(978)
		x =             -290; #20833; // Sample(979)
		x =             -183; #20833; // Sample(980)
		x =                0; #20833; // Sample(981)
		x =              183; #20833; // Sample(982)
		x =              290; #20833; // Sample(983)
		x =              277; #20833; // Sample(984)
		x =              150; #20833; // Sample(985)
		x =              -39; #20833; // Sample(986)
		x =             -212; #20833; // Sample(987)
		x =             -297; #20833; // Sample(988)
		x =             -260; #20833; // Sample(989)
		x =             -115; #20833; // Sample(990)
		x =               78; #20833; // Sample(991)
		x =              238; #20833; // Sample(992)
		x =              300; #20833; // Sample(993)
		x =              238; #20833; // Sample(994)
		x =               78; #20833; // Sample(995)
		x =             -115; #20833; // Sample(996)
		x =             -260; #20833; // Sample(997)
		x =             -297; #20833; // Sample(998)
		x =             -212; #20833; // Sample(999)
		x =              -39; #20833; // Sample(1000)
        $stop;
    end
endmodule
